* -- Netlist template

* --- Voltage Sources ---

Vd Vd 0 0

Vg Vg 0 0

Vs Vs 0 0

Vb Vb 0 0


* --- Transistor ---
mbsim4  Vd  Vg  Vs  Vb  nmos  AD=0.194e-12  AS=0.194e-12  NF=1  W=3.60E-07  L=1.80E-07  RGEOMOD=0  PD=1.8e-6  PS=1.8E-6 
.MODEL nmos nmos  WMAX=1  WMIN=0  LMAX=1  LMIN=0  WWLC=0  WLC=0  WLC=0  LWLC=0  LWC=0  LLC=0  LWL=0  LWN=1  LW=0  LLN=1  LL=0  WWL=0  WWN=1  WW=0  WLN=1  WL=0  NJD=1  NJd=1  TCJSWG=0  TCJSW=0  TCJ=0  TPBSWG=0  TPBSW=0  TPB=0  XTIS=3  NJS=1  PRT=0  AT=3.30E+04  UC1=0.025  UB1=-1.00E-18  UA1=1.00E-09  KT2=0.022  KT1L=0  KT1=-0.11  UTE=-1.5  TNOM=27  XTID=3  XTID=3  PBSWGD=1  PBSWGS=1  PBSWD=1  PBSWS=1  PBS=1  PBD=1  MJSWGD=0.33  MJSWGS=0.33  CJSWGD=5.00E-10  CJSWGS=5.00E-10  CJSWD=5.00E-10  CJSWS=5.00E-10  MJSWD=0.33  MJSWS=0.33  MJD=0.5  MJS=0.5  CJD=5.00E-04  CJS=5.00E-04  JSWGD=0  JSWGS=0  JSWD=0  JSWS=0  JSD=1.00E-04  JSS=1.00E-04  BVD=10  BVS=10  XJBVD=1  XJBVS=1  IJTHDFWD=0.1  IJTHSFWD=0.1  IJTHDREV=0.1  IJTHSREV=0.1  NGCON=1  XGL=0  XGW=0  MIN=0  DWJ=0  DMCGT=0  DMDG=0  DMCI=0  DMCG=0  TNOIB=3.5  TNOIA=1.5  NTNOI=1  KF=0  EF=1  AF=1  EM=4.10E+07  NOIC=8.75  NOIB=3.125e26  NOIA=6.25e41  GBMIN=1.00E-12  RBSB=50  RBDB=50  RBPS=50  RBPD=50  RBPB=50  XRCRG2=1  XRCRG1=12  MOIN=15  ACDE=1  VOFFCV=0  NOFF=1  VFBCV=-1  DWC=0  DLC=0  CLE=0.6  CLC=1.00E-07  CF=0  CKAPPAD=0.6  CKAPPAS=0.6  CGDL=0  CGSL=0  CGBO=0  CGDO=0  CGSO=0  XPART=0  TOXREF=3.00E-09  NTOX=1  PIGCD=1  POXEDGE=1  NIGC=1  DLCIG=0  CIGSD=0.075  BIGSD=0.054  AIGSD=0.43  CIGC=0.075  BIGC=0.054  AIGC=0.054  NIGBINV=3  EIGBINV=1.1  CIGBINV=0.006  BIGBINV=0.03  AIGBINV=0.35  NIGBACC=1  CIGBACC=0.075  BIGBACC=0.054  AIGBACC=0.43  DGIDL=0.8  CGIDL=0.5  BGIDL=2.30E+09  AGIDL=0  BETA0=30  ALPHA1=0  ALPHA0=0  NRD=1  NRS=1  WR=1  PRWB=0  PRWG=1  RSWMIN=0  RSW=100  RDWMIN=0  RDW=100  RDSWMIN=0  RDSW=200  PDITSD=0  PDITSL=0  PDITS=0  FPROUT=0  DELTA=0.01  PVAG=0  PSCBE2=1.00E-05  PSCBE1=4.24E+08  DROUT=0.56  PDIBLCB=0  PDIBLC2=0.0086  PDIBLC1=0.39  PCLM=1.3  CDSCD=0  CDSCB=0  CDSC=2.40E-04  CIT=0  DSUB=0.56  ETAB=-0.07  ETA0=0.08  NFACTOR=1  MINV=0  VOFFL=0  VOFF=-0.08  DWB=0  DWG=0  LINT=0  WINT=0  A2=1  A1=0  KETA=-0.047  B1=0  B0=0  AGS=0  A0=1  VSAT=8.00E+04  EU=1.67  UC=-0.0465  UB=1.00E-19  UA=1.0e-9  U0=0.067  DVT2W=-0.032  DVT1W=5.30E+06  DVT0W=0  DVTP1=0  DVTP0=0  DVT2=-0.032  DVT1=0.53  DVT0=2.2  VBM=-3  LPEB=0  LPE0=1.74E-07  W0=2.50E-06  K3B=0  K3=80  K2=0  K1=0.5  PHIN=0  VFB=-1  VTH0=0.7  RSHG=0.1  RSH=0  XT=1.55E-07  NSD=1.00E+20  NGATE=0  NSUB=6.00E+16  NDEP=1.70E+17  XJ=1.50E-07  DTOX=0  TOXM=3.0E-9  TOXP=3e-9  TOXE=3.00E-09  EPSROX=3.9  TYPE=1  GEOMOD=0  PERMOD=1  DIOMOD=1  TNOIMOD=0  FNOIMOD=1  ACNQSMOD=0  TRNQSMOD=0  RBODYMOD=0  RGATEMOD=0  CAPMOD=2  IGBMOD=0  IGCMOD=0  RDSMOD=0  MOBMOD=1  PARAMCHK=1  BINUNIT=1  VERSION=4.0  LEVEL=14 

* --- Transfer ---
.control

save all
save  i(vs) i(vd) i(vg) i(vb) @mbsim4[qd] @mbsim4[qg] @mbsim4[qb] @mbsim4[cdd] @mbsim4[cdg] @mbsim4[cds] @mbsim4[cgd] @mbsim4[cgg] @mbsim4[cgs] @mbsim4[cbd] @mbsim4[cbg] @mbsim4[cbs] @mbsim4[gm] @mbsim4[gds] 

dc  Vd 0 1 0.1  Vg 0 1 0.1 

wrdata output  i(vs) i(vd) i(vg) i(vb) @mbsim4[qd] @mbsim4[qg] @mbsim4[qb] @mbsim4[cdd] @mbsim4[cdg] @mbsim4[cds] @mbsim4[cgd] @mbsim4[cgg] @mbsim4[cgs] @mbsim4[cbd] @mbsim4[cbg] @mbsim4[cbs] @mbsim4[gm] @mbsim4[gds] 

.endc

.end